library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fsm is
	port(en,reset_n,clk,config,ini_pausa,jugador_act,min_value_j0,min_value_j1,mov_j0_gt40,mov_j1_gt40: in std_logic;
																		modo: in std_logic_vector(1 downto 0);
									ini_pausa_j0,borrar_j0,ini_pausa_j1,borrar_j1,en_sel,en_j1,en_j0:out std_logic);
end fsm;

architecture arch of fsm is
	type estados is (ST_IDLE,ST_WAIT_CONFIG,ST_PLAYERS_CONFIG, ST_PLAYER_0_P,ST_PLAYER_1_P,ST_PLAYER_0,ST_PLAYER_1,ST_PLAYER_0_L,ST_PLAYER_1_L,ST_PLAYER_0_M,ST_PLAYER_1_M);
	signal state_reg, state_next: estados;
	begin
		process(reset_n,en,clk)
			begin
				if reset_n = '0' then
					state_reg <= ST_IDLE;
				elsif rising_edge(clk) then
					if (en='1') then
						state_reg <= state_next;
					else
						state_reg <= state_reg;
					end if;
				end if;
		end process;
		
		process(state_reg,config,ini_pausa,jugador_act,min_value_j0,min_value_j1,reset_n)
			begin
				case state_reg is
					when ST_IDLE =>
						if config = '0' then
							state_next <= ST_IDLE;
						elsif config = '1' then
							state_next <= ST_WAIT_CONFIG;
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '1';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '1';
						
					when ST_WAIT_CONFIG =>
						if config = '1' then
							state_next <= ST_WAIT_CONFIG;
						elsif config ='0' then
							state_next <= ST_PLAYERS_CONFIG;
						end if;
						en_sel <= '1';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '1';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '1';	
						
					when ST_PLAYERS_CONFIG =>
						if ini_pausa='1' then
							if jugador_act = '1' then
								state_next <= ST_PLAYER_1_P;
							elsif jugador_act = '0' then
								state_next <= ST_PLAYER_0_P;
							end if;
						else
							state_next <= ST_PLAYERS_CONFIG;
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
					when ST_PLAYER_0_P =>
						if ini_pausa = '1' then
							state_next <= ST_PLAYER_0;
						else
							state_next <= ST_PLAYER_0_P;
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';			
						
					when ST_PLAYER_1_P =>
						if ini_pausa = '1' then
							state_next <= ST_PLAYER_1;
						else
							state_next <= ST_PLAYER_1_P;
						end if;				
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
					when ST_PLAYER_0 =>
						if ini_pausa = '0' then
							state_next <= ST_PLAYER_0_P;
						elsif min_value_j0 = '1' then
							state_next <= ST_PLAYER_0_L;
						elsif jugador_act = '1' then
							state_next <= ST_PLAYER_0_M;---cambiado
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '1';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
					when ST_PLAYER_1 => 
						if ini_pausa = '0' then
							state_next <= ST_PLAYER_1_P;
						elsif min_value_j1 = '1' then
							state_next <= ST_PLAYER_1_L;
						elsif jugador_act = '0' then
							state_next <= ST_PLAYER_1_M;--cambiado
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '1';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
					when ST_PLAYER_1_M =>
						state_next <= ST_PLAYER_0;
 						en_sel <= '0';
						en_j1 <= '1';--añadido
						ini_pausa_j0 <= '1';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';

					when ST_PLAYER_0_M =>
						state_next <= ST_PLAYER_1;
 						en_sel <= '0';
						en_j0 <= '1';--añadido
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '1';
						borrar_j1 <= '0';						
						
					when ST_PLAYER_0_L =>
						if reset_n = '0'then
							state_next <= ST_IDLE;
						else
							state_next <= ST_PLAYER_0_L;
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
					when ST_PLAYER_1_L =>
						if reset_n = '0' then
							state_next <= ST_IDLE;
						else
							state_next <= ST_PLAYER_1_L;
						end if;
						en_sel <= '0';
						ini_pausa_j0 <= '0';
						borrar_j0 <= '0';
						ini_pausa_j1 <= '0';
						borrar_j1 <= '0';
						en_j0 <= '0';
						en_j1 <= '0';
						
				end case;
		end process;
end arch;